module timer(
    
);
    
endmodule