module FIFO #(parameter FIFO_WIDTH = 9)
(
    input clk,rst_n,wr_en,rd_en,
    input [FIFO_WIDTH-1:0]data_in,
    output full,almostfull,empty,almostempty,
    output reg overflow,underflow,
    output reg [FIFO_WIDTH-1:0]data_out,
    output reg wr_ack
);

parameter FIFO_DEPTH = 16;
localparam max_fifo_addr = $clog2(FIFO_DEPTH);
reg [FIFO_WIDTH-1:0]mem[FIFO_DEPTH-1:0];
reg [max_fifo_addr-1:0] wr_ptr, rd_ptr;
reg [max_fifo_addr:0] count;

always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        wr_ptr <= 0;
		wr_ack <= 0;
		overflow <= 0;
    end
    else if (wr_en && count < FIFO_DEPTH) begin
        mem[wr_ptr] <= data_in;
        wr_ack <= 1;
        wr_ptr <= wr_ptr + 1;
        overflow <= 0;
    end
    else begin
        wr_ack <= 0;
        if(wr_en && full) begin
            overflow <= 1;
        end
        else begin
            overflow <= 0;
        end
    end
end

always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        rd_ptr <= 0;
		underflow <= 0;
    end
    else if (rd_en && count > 0) begin
        data_out <= mem[rd_ptr];
        rd_ptr <= rd_ptr + 1;
        underflow <= 0;
    end
    else begin
        if(empty && rd_en) begin
			underflow <= 1;
		end
		else begin
			underflow <= 0;
		end
    end
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n) begin
		count <= 0;
	end
	else begin
		if	((({wr_en, rd_en} == 2'b10) && !full)) 
			count <= count + 1;
		else if ((({wr_en, rd_en} == 2'b01) && !empty))
			count <= count - 1;
			else if(({wr_en, rd_en} == 2'b11)) begin 
				if(full)
				count <= count - 1;
				else if(empty)
				count <= count + 1;
			end
	end
end

assign full = (count == FIFO_DEPTH)? 1 : 0;
assign empty = (count == 0)? 1 : 0;
assign almostfull = (count == FIFO_DEPTH-1)? 1 : 0; 
assign almostempty = (count == 1)? 1 : 0;
endmodule